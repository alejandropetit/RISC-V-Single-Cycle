module control #(parameter XLEN=32)(input logic clk, reset, SrcBCtrl, input logic [XLEN-1:0] PC, Instr, output logic [3:0] AluCtrl, output logic [1:0] ExtCtrl);

endmodule